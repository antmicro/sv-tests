// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: net_decl_assignment
:description: net declaration assignment test
:tags: 10.3.1
:results_group: ten-three
*/
module top(input a, input b);

wire w = a & b;

endmodule
